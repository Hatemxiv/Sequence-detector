// Copyright (C) 2022  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 22.1std.0 Build 915 10/25/2022 SC Standard Edition
// Created on Sat Nov  4 18:48:45 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    reset,clock,serial_in,start,
    seq_out);

    input reset;
    input clock,start;
    input serial_in;
    tri0 reset;
    tri0 serial_in;
    output seq_out;
    reg seq_out;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter s0=0,s1=1,s2=2,s3=3,s4=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or serial_in)
    begin
        if (reset) begin
            reg_fstate <= s0;
            seq_out <= 1'b0;
        end
        else if(start) begin
            seq_out <= 1'b0;
            case (fstate)
                s0: begin
                    if ((serial_in == 1'b1))
                        reg_fstate <= s1;
                    else if ((serial_in == 1'b0))
                        reg_fstate <= s0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s0;

                    seq_out <= 1'b0;
                end
                s1: begin
                    if ((serial_in == 1'b0))
                        reg_fstate <= s2;
                    else if ((serial_in == 1'b1))
                        reg_fstate <= s1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s1;

                    seq_out <= 1'b0;
                end
                s2: begin
                    if ((serial_in == 1'b0))
                        reg_fstate <= s0;
                    else if ((serial_in == 1'b1))
                        reg_fstate <= s3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s2;

                    seq_out <= 1'b0;
                end
                s3: begin
                    if ((serial_in == 1'b1))
                        reg_fstate <= s4;
                    else if ((serial_in == 1'b0))
                        reg_fstate <= s2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s3;

                    seq_out <= 1'b0;
                end
                s4: begin
                    if ((serial_in == 1'b0))
                        reg_fstate <= s0;
                    else if ((serial_in == 1'b1))
                        reg_fstate <= s1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s4;

                    seq_out <= 1'b1;
                end
                default: begin
                    seq_out <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
